module counter();

endmodule
